*id vs vds
.include ALD1105.txt
m1 1 2 0 4 ALD1105P 
vgs 2 0 -5
vd 1 3 0V
vsb 4 0 4
vds 3 0 200m
.control
dc vgs 0 -5 -0.02 vsb 0 4 1
plot i(vd)
hardcopy p1 i(vd)
wrdata p1_data i(vd)
.endc
.end 


