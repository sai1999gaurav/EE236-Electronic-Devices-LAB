*id vs vds
.include ALD1107.txt
m1 1 2 0 0 ALD1107 
vgs 0 2 1.5V
vd 1 3 0V
vds 3 0 -5
.control
dc vds 0 -5 -0.02 vgs 1.5 3 0.5
plot -i(vd) 
hardcopy p1 -i(vd)
wrdata p1_data -i(vd)
.endc
.end 


